`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:03:12 03/08/2020 
// Design Name: 
// Module Name:    Left_shifter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: [ 
//
//////////////////////////////////////////////////////////////////////////////////
module Left_shifter( input [31:0]a, input [4:0]b, output [31:0]c);
wire [31:0]w0;
wire [31:0]w1;
wire [31:0]w2;
wire [31:0]w3;

mux_8_chain stage0(.in0(a), .out(w0), .Select(b[0]),
						.in1({a[30], a[29], a[28], a[27], a[26], a[25], a[24], a[23], 
						       a[22], a[21], a[20], a[19], a[18], a[17], a[16], a[15],
								 a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7],
								 a[6], a[5], a[4], a[3], a[2], a[1], a[0], a[31]})
);

mux_8_chain stage1(.in0(w0), .out(w1), .Select(b[1]),
                   .in1({w0[29], w0[28], w0[27], w0[26], w0[25], w0[24], w0[23], w0[22], 
						       w0[21], w0[20], w0[19], w0[18], w0[17], w0[16], w0[15], w0[14],
								 w0[13], w0[12], w0[11], w0[10], w0[9], w0[8], w0[7], w0[6],
								 w0[5], w0[4], w0[3], w0[2], w0[1], w0[0], w0[31], w0[30]})
);

mux_8_chain stage2(.in0(w1), .out(w2), .Select(b[2]),
                   .in1({w1[27], w1[26], w1[25], w1[24], w1[23], w1[22], w1[21], w1[20], 
						       w1[19], w1[18], w1[17], w1[16], w1[15], w1[14], w1[13], w1[12],
								 w1[11], w1[10], w1[9], w1[8], w1[7], w1[6], w1[5], w1[4],
								 w1[3], w1[2], w1[1], w1[0], w1[31], w1[30], w1[29], w1[28]})
);

mux_8_chain stage3(.in0(w2), .out(w3), .Select(b[3]),
                   .in1({w2[23], w2[22], w2[21], w2[20], w2[19], w2[18], w2[17], w2[16], 
						       w2[15], w2[14], w2[13], w2[12], w2[11], w2[10], w2[9], w2[8],
								 w2[7], w2[6], w2[5], w2[4], w2[3], w2[2], w2[1], w2[0],
								 w2[31], w2[30], w2[29], w2[28], w2[27], w2[26], w2[25], w2[24]})
);

mux_8_chain stage4(.in0(w3), .out(c), .Select(b[4]),
                   .in1({w3[15], w3[14], w3[13], w3[12], w3[11], w3[10], w3[9], w3[8], 
						       w3[7], w3[6], w3[5], w3[4], w3[3], w3[2], w3[1], w3[0],
								 w3[31], w3[30], w3[29], w3[28], w3[27], w3[26], w3[25], w3[24],
								 w3[23], w3[22], w3[21], w3[20], w3[19], w3[18], w3[17], w3[16]})
	
);

endmodule
